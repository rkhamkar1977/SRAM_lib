module decoder_2( address_1,
                  address_2,
                  read_enable,
                  write_enable,
                  read_wl1,
                  read_wl2,
                  write_wl
                );

    input       [6:0]   address_1;
    input       [6:0]   address_2;
    input       [1:0]   read_enable;
    input               write_enable;
    output  reg [127:0] read_wl1;
    output  reg [127:0] read_wl2;
    output  reg [127:0] write_wl;

    
    always @(*) begin
        case (address_1)
            7'd0: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001 : 0;
            end
            7'd1: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010 : 0;
            end
            7'd2: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100 : 0;
            end
            7'd3: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000 : 0;
            end
            7'd4: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000 : 0;
            end
            7'd5: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000 : 0;
            end
            7'd6: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000 : 0;
            end
            7'd7: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000 : 0;
            end
            7'd8: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000 : 0;
            end
            7'd9: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000 : 0;
            end
            7'd10: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000 : 0;
            end
            7'd11: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000 : 0;
            end
            7'd12: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000 : 0;
            end
            7'd13: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000 : 0;
            end
            7'd14: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000 : 0;
            end
            7'd15: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000 : 0;
            end
            7'd16: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000 : 0;
            end
            7'd17: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000 : 0;
            end
            7'd18: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000 : 0;
            end
            7'd19: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000 : 0;
            end
            7'd20: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000 : 0;
            end
            7'd21: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000 : 0;
            end
            7'd22: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000 : 0;
            end
            7'd23: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000 : 0;
            end
            7'd24: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000 : 0;
            end
            7'd25: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000 : 0;
            end
            7'd26: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000 : 0;
            end
            7'd27: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000 : 0;
            end
            7'd28: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000 : 0;
            end
            7'd29: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000 : 0;
            end
            7'd30: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000 : 0;
            end
            7'd31: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000 : 0;
            end
            7'd32: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000 : 0;
            end
            7'd33: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000 : 0;
            end
            7'd34: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000 : 0;
            end
            7'd35: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000 : 0;
            end
            7'd36: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000 : 0;
            end
            7'd37: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000 : 0;
            end
            7'd38: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000 : 0;
            end
            7'd39: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000 : 0;
            end
            7'd40: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000 : 0;
            end
            7'd41: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000 : 0;
            end
            7'd42: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000 : 0;
            end
            7'd43: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000 : 0;
            end
            7'd44: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000 : 0;
            end
            7'd45: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000 : 0;
            end
            7'd46: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000 : 0;
            end
            7'd47: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000 : 0;
            end
            7'd48: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000 : 0;
            end
            7'd49: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000 : 0;
            end
            7'd50: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000 : 0;
            end
            7'd51: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd52: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd53: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd54: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd55: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd56: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd57: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd58: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd59: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd60: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd61: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd62: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd63: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd64: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd65: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd66: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd67: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd68: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd69: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd70: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd71: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd72: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd73: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd74: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd75: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd76: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd77: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd78: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd79: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd80: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd81: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd82: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd83: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd84: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd85: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd86: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd87: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd88: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd89: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd90: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd91: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd92: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd93: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd94: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd95: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd96: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd97: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd98: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd99: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd100: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd101: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd102: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd103: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd104: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd105: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd106: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd107: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd108: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd109: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd110: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd111: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd112: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd113: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd114: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd115: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd116: begin 
                read_wl1 = read_enable[0] ? 128'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd117: begin 
                read_wl1 = read_enable[0] ? 128'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd118: begin 
                read_wl1 = read_enable[0] ? 128'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd119: begin 
                read_wl1 = read_enable[0] ? 128'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd120: begin 
                read_wl1 = read_enable[0] ? 128'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd121: begin 
                read_wl1 = read_enable[0] ? 128'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd122: begin 
                read_wl1 = read_enable[0] ? 128'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd123: begin 
                read_wl1 = read_enable[0] ? 128'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd124: begin 
                read_wl1 = read_enable[0] ? 128'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd125: begin 
                read_wl1 = read_enable[0] ? 128'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd126: begin 
                read_wl1 = read_enable[0] ? 128'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd127: begin 
                read_wl1 = read_enable[0] ? 128'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
                write_wl = write_enable ? 128'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
        endcase
        case (address_2) 
            7'd0: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001 : 0;
            end
            7'd1: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010 : 0;
            end
            7'd2: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100 : 0;
            end
            7'd3: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000 : 0;
            end
            7'd4: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000 : 0;
            end
            7'd5: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000 : 0;
            end
            7'd6: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000 : 0;
            end
            7'd7: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000 : 0;
            end
            7'd8: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000 : 0;
            end
            7'd9: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000 : 0;
            end
            7'd10: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000 : 0;
            end
            7'd11: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000 : 0;
            end
            7'd12: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000 : 0;
            end
            7'd13: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000 : 0;
            end
            7'd14: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000 : 0;
            end
            7'd15: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000 : 0;
            end
            7'd16: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000 : 0;
            end
            7'd17: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000 : 0;
            end
            7'd18: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000 : 0;
            end
            7'd19: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000 : 0;
            end
            7'd20: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000 : 0;
            end
            7'd21: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000 : 0;
            end
            7'd22: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000 : 0;
            end
            7'd23: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000 : 0;
            end
            7'd24: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000 : 0;
            end
            7'd25: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000 : 0;
            end
            7'd26: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000 : 0;
            end
            7'd27: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000 : 0;
            end
            7'd28: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000 : 0;
            end
            7'd29: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000 : 0;
            end
            7'd30: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000 : 0;
            end
            7'd31: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000 : 0;
            end
            7'd32: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000 : 0;
            end
            7'd33: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000 : 0;
            end
            7'd34: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000 : 0;
            end
            7'd35: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000 : 0;
            end
            7'd36: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000 : 0;
            end
            7'd37: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000 : 0;
            end
            7'd38: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000 : 0;
            end
            7'd39: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000 : 0;
            end
            7'd40: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000 : 0;
            end
            7'd41: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000 : 0;
            end
            7'd42: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000 : 0;
            end
            7'd43: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000 : 0;
            end
            7'd44: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000 : 0;
            end
            7'd45: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000 : 0;
            end
            7'd46: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000 : 0;
            end
            7'd47: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000 : 0;
            end
            7'd48: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000 : 0;
            end
            7'd49: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000 : 0;
            end
            7'd50: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000 : 0;
            end
            7'd51: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd52: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd53: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd54: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd55: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd56: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd57: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd58: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd59: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd60: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd61: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd62: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd63: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd64: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd65: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd66: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd67: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd68: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd69: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd70: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd71: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd72: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd73: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd74: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd75: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd76: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd77: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd78: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd79: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd80: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd81: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd82: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd83: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd84: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd85: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd86: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd87: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd88: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd89: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd90: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd91: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd92: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd93: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd94: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd95: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd96: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd97: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd98: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd99: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd100: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd101: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd102: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd103: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd104: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd105: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd106: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd107: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd108: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd109: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd110: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd111: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd112: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd113: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd114: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd115: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd116: begin 
                read_wl2 = read_enable[1] ? 128'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd117: begin 
                read_wl2 = read_enable[1] ? 128'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd118: begin 
                read_wl2 = read_enable[1] ? 128'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd119: begin 
                read_wl2 = read_enable[1] ? 128'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd120: begin 
                read_wl2 = read_enable[1] ? 128'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd121: begin 
                read_wl2 = read_enable[1] ? 128'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd122: begin 
                read_wl2 = read_enable[1] ? 128'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd123: begin 
                read_wl2 = read_enable[1] ? 128'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd124: begin 
                read_wl2 = read_enable[1] ? 128'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd125: begin 
                read_wl2 = read_enable[1] ? 128'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd126: begin 
                read_wl2 = read_enable[1] ? 128'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
            7'd127: begin 
                read_wl2 = read_enable[1] ? 128'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : 0;
            end
        endcase
    end

endmodule
